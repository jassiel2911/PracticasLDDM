library verilog;
use verilog.vl_types.all;
entity Segunda_Parte_vlg_vec_tst is
end Segunda_Parte_vlg_vec_tst;
