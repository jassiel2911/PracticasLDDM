library verilog;
use verilog.vl_types.all;
entity Segunda_Parte_vlg_check_tst is
    port(
        X               : in     vl_logic;
        Y               : in     vl_logic;
        Z               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Segunda_Parte_vlg_check_tst;
