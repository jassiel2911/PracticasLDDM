library verilog;
use verilog.vl_types.all;
entity Ejercicio_Previo_vlg_vec_tst is
end Ejercicio_Previo_vlg_vec_tst;
