library verilog;
use verilog.vl_types.all;
entity anodo_vlg_vec_tst is
end anodo_vlg_vec_tst;
