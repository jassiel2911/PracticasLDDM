library verilog;
use verilog.vl_types.all;
entity codvhd1_vlg_check_tst is
    port(
        P               : in     vl_logic;
        S               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end codvhd1_vlg_check_tst;
