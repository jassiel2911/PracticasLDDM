library verilog;
use verilog.vl_types.all;
entity codvhd1_vlg_vec_tst is
end codvhd1_vlg_vec_tst;
